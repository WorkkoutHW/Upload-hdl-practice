module GATE_AND(input A, B, C);

assign C = A & B;

endmodule